// ============================================================
// itch_reset.vh
// Universal reset logic macro, delegates to decoder-specific field resets
// ============================================================

`define ITCH_RESET_LOGIC \
    `ITCH_RESET_FIELDS
